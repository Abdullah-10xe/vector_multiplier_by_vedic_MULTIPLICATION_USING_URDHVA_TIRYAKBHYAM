module  multiplier_16bit  (input  logic clk, input logic rst,
                           input  logic [15:0] operand_a_16bit,
                           input  logic [15:0] operand_b_16bit,
                           input  logic [1:0] precision,
                           output logic [31:0] output_16bit_mul);
  logic [3:0][15:0]in_8bit_mul_block;
  logic [31:0]     output_16bit_mul_wire; 
  logic [31:0] output_16bit_mul_pr8;
  logic [31:0] output_16bit_mul_pr16;
  logic [7:0]  mux_a_8bit_pre;
  logic [15:0] csa_sum;
  logic [15:0] csa_carry;
  logic        carry_bka;
  logic        mux_sel;
 
  
  multiplier_8bit unit2_0 (.operand_a_8bit(operand_a_16bit[7:0]),.operand_b_8bit(operand_b_16bit[7:0]),.output_8bit_mul(in_8bit_mul_block[0]));
  multiplier_8bit unit2_1 (.operand_a_8bit(mux_a_8bit_pre),.operand_b_8bit( operand_b_16bit[15:8]),.output_8bit_mul(in_8bit_mul_block[1]));
  multiplier_8bit unit2_2 (.operand_a_8bit(operand_a_16bit[15:8]),.operand_b_8bit(operand_b_16bit[7:0]),.output_8bit_mul(in_8bit_mul_block[2]));
  multiplier_8bit unit2_3 (.operand_a_8bit(operand_a_16bit[15:8]),.operand_b_8bit(operand_b_16bit[15:8]),.output_8bit_mul(in_8bit_mul_block[3]));
  
  
  
  carry_save_adder #(.ADDER_WIDTH(16)) cs_adder (
    .operand_a_csa({in_8bit_mul_block [3][7:0],in_8bit_mul_block [0][15:8]}), 
    .operand_b_csa(in_8bit_mul_block[1]),
    .operand_c_csa(in_8bit_mul_block[2]),
    .sum_csv(csa_sum),
    .carry_csv(csa_carry)
    );
  
  
  
  brent_kung_adder #(.ADDER_WIDTH(16),.NO_CARRY(0)) bk_adder  (
    .operand_a_bka({in_8bit_mul_block[3][8], csa_sum[15:1]}), 
    .operand_b_bka(csa_carry),                     
    .sum_bka(output_16bit_mul_pr16[24:9]),
     .carry_bka(carry_bka)
);
  
  carray_select_adder #(.ADDER_WIDTH(7)) csela (  
                                        .operand_a_csela(in_8bit_mul_block[3][15:9]),
                                       .carry_in_csela(carry_bka),
                                       .sum_csela(output_16bit_mul_pr16[31:25]));
     
  
  
  
  assign mux_sel=(precision==2'b00);
  assign output_16bit_mul_pr16 [8:0]={csa_sum[0],in_8bit_mul_block[0][7:0]};
  assign output_16bit_mul_pr8 ={in_8bit_mul_block[1],in_8bit_mul_block[0]};
  assign mux_a_8bit_pre=mux_sel?operand_a_16bit[15:8]:operand_a_16bit[7:0];
  assign output_16bit_mul_wire=mux_sel?output_16bit_mul_pr8 :output_16bit_mul_pr16  ;

  
  
  always_ff @(posedge clk,negedge rst)
    begin
      if(!rst)
        begin
         output_16bit_mul<=0;
        
        end
        else
          begin
          
      output_16bit_mul=output_16bit_mul_wire;
     
          end
      end
    
    
      
    
    
    
 
endmodule


